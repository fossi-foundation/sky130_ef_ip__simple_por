magic
tech sky130A
magscale 1 2
timestamp 1747235245
<< isosubstrate >>
rect 1330 7236 8715 11911
rect 234 0 8715 7236
<< nwell >>
rect 1383 7415 1885 10884
rect 889 84 1340 6666
<< pwell >>
rect 2658 2649 2868 2867
rect 2105 477 2115 533
<< psubdiff >>
rect 44 11784 116 11808
rect 44 52 116 76
<< mvpsubdiff >>
rect 8319 10986 8648 11020
rect 1229 7452 1297 10870
rect 1956 7004 2358 7028
rect 1956 3178 2358 3202
<< mvnsubdiff >>
rect 1449 7481 1483 10841
<< psubdiffcont >>
rect 44 76 116 11784
<< mvpsubdiffcont >>
rect 1956 3202 2358 7004
<< locali >>
rect 8 11792 132 11832
rect 1362 11817 8638 11872
rect 1362 10883 1386 11817
rect 1437 11800 8638 11817
rect 1437 10883 1483 11800
rect 1534 10894 8648 11020
rect 1362 10840 1483 10883
rect 2263 10870 8648 10894
rect 2263 10840 2541 10870
rect 1362 7481 1449 10840
rect 1362 7148 1483 7481
rect 2297 7148 2541 10840
rect 2655 10670 2871 10851
rect 8303 10669 8519 10849
rect 2655 9512 2871 9899
rect 8303 9897 8519 10284
rect 2655 8740 2871 9127
rect 8303 9125 8519 9512
rect 2655 7968 2871 8355
rect 8303 8353 8519 8740
rect 2655 7196 2871 7583
rect 8303 7581 8519 7968
rect 398 7131 1679 7148
rect 398 6950 411 7131
rect 572 7124 1679 7131
rect 572 6950 1249 7124
rect 398 6941 1249 6950
rect 1662 6941 1679 7124
rect 398 6905 1679 6941
rect 1229 3057 1679 6905
rect 1846 7004 2541 7148
rect 1846 3202 1956 7004
rect 2358 6130 2541 7004
rect 2655 6424 2871 6811
rect 8303 6809 8519 7196
rect 2431 3234 2541 6130
rect 2655 5652 2871 6039
rect 8303 6037 8519 6424
rect 2655 4880 2871 5267
rect 8303 5265 8519 5652
rect 2655 4108 2871 4495
rect 8303 4493 8519 4880
rect 2655 3336 2871 3723
rect 8303 3721 8519 4108
rect 2358 3202 2541 3234
rect 1233 197 1379 3057
rect 1846 2965 2541 3202
rect 1846 2921 2364 2965
rect 396 183 1379 197
rect 396 71 409 183
rect 494 71 1379 183
rect 2296 519 2364 2921
rect 2493 703 2541 2965
rect 2655 2854 2871 2951
rect 8303 2949 8519 3336
rect 2655 2662 2669 2854
rect 2855 2662 2871 2854
rect 2655 2564 2871 2662
rect 2655 1792 2871 2179
rect 8303 2177 8519 2564
rect 2655 1020 2871 1407
rect 8303 1405 8519 1792
rect 2493 519 2871 703
rect 8303 633 8519 1020
rect 2296 300 2871 519
rect 2296 135 2366 300
rect 396 55 1379 71
rect 1505 62 2366 135
rect 2492 62 2871 300
rect 8303 65 8519 248
rect 1505 49 2871 62
rect 8 0 132 40
<< viali >>
rect 8 11784 132 11792
rect 8 76 44 11784
rect 44 76 116 11784
rect 116 76 132 11784
rect 1386 10883 1437 11817
rect 1814 11323 2405 11363
rect 805 10799 1001 10833
rect 883 9473 930 9810
rect 624 9238 830 9284
rect 883 7618 930 7821
rect 1788 10284 1949 10330
rect 1917 8664 1964 8867
rect 1806 8453 2000 8520
rect 1850 7884 1909 8142
rect 2654 10216 3086 10354
rect 411 6950 572 7131
rect 1249 6941 1662 7124
rect 1991 3234 2358 6130
rect 2358 3234 2431 6130
rect 8 40 132 76
rect 409 71 494 183
rect 2364 519 2493 2965
rect 2669 2662 2855 2854
rect 2366 62 2492 300
<< metal1 >>
rect 0 11792 140 11832
rect 0 40 8 11792
rect 132 40 140 11792
rect 1360 11817 8638 11840
rect 406 10816 559 11624
rect 956 10919 1010 10929
rect 406 7332 432 10816
rect 531 7332 559 10816
rect 793 10833 956 10839
rect 793 10799 805 10833
rect 793 10793 956 10799
rect 1010 10793 1013 10839
rect 956 10757 1010 10767
rect 1114 10663 1267 11619
rect 631 10304 685 10314
rect 631 10142 685 10152
rect 633 9290 683 10142
rect 877 9810 936 9822
rect 877 9473 883 9810
rect 930 9473 936 9810
rect 612 9284 842 9290
rect 612 9238 624 9284
rect 830 9238 842 9284
rect 612 9232 842 9238
rect 877 8533 936 9473
rect 877 7821 936 8353
rect 877 7618 883 7821
rect 930 7618 936 7821
rect 877 7606 936 7618
rect 1114 8632 1141 10663
rect 1235 8632 1267 10663
rect 1114 8357 1267 8632
rect 406 7298 559 7332
rect 1114 7320 1141 8357
rect 1235 7320 1267 8357
rect 1114 7293 1267 7320
rect 1360 10883 1386 11817
rect 1437 11802 8638 11817
rect 1556 11731 1608 11802
rect 4718 11731 5004 11802
rect 8605 11731 8638 11802
rect 1556 11692 8638 11731
rect 1556 11256 1591 11692
rect 2619 11566 8453 11591
rect 2619 11550 4950 11566
rect 2619 11482 2645 11550
rect 4893 11498 4950 11550
rect 8431 11498 8453 11566
rect 4893 11482 5066 11498
rect 2619 11460 5066 11482
rect 6165 11481 8453 11498
rect 1782 11379 2440 11386
rect 1782 11310 1797 11379
rect 2413 11310 2440 11379
rect 1782 11304 2440 11310
rect 1437 11227 1591 11256
rect 1437 10883 1482 11227
rect 1533 11105 8670 11128
rect 1533 11031 2014 11105
rect 8634 11031 8670 11105
rect 1533 10980 8670 11031
rect 1360 10846 1482 10883
rect 2153 10923 2365 10980
rect 1360 10764 1591 10846
rect 1360 8616 1385 10764
rect 1560 10530 1591 10764
rect 1850 10686 1919 10696
rect 1560 8616 1590 10530
rect 1850 10336 1919 10521
rect 2153 10545 2177 10923
rect 2248 10545 2365 10923
rect 2605 10819 8673 10881
rect 1776 10330 1961 10336
rect 1776 10284 1788 10330
rect 1949 10284 1961 10330
rect 1776 10278 1961 10284
rect 2153 10082 2365 10545
rect 2414 10714 2508 10730
rect 2414 10247 2424 10714
rect 2497 10329 2508 10714
rect 2639 10354 3102 10367
rect 2639 10329 2654 10354
rect 2497 10247 2654 10329
rect 2414 10235 2654 10247
rect 2639 10216 2654 10235
rect 3086 10216 3102 10354
rect 2639 10201 3102 10216
rect 1360 8334 1590 8616
rect 1911 8867 1970 8879
rect 1911 8664 1917 8867
rect 1964 8664 1970 8867
rect 1911 8530 1970 8664
rect 1806 8526 2000 8530
rect 1794 8520 2012 8526
rect 1794 8453 1806 8520
rect 2000 8453 2012 8520
rect 1794 8447 2012 8453
rect 1806 8443 2000 8447
rect 1360 7185 1385 8334
rect 1560 7185 1590 8334
rect 1360 7148 1590 7185
rect 1844 8142 1915 8154
rect 1844 7884 1850 8142
rect 1909 7884 1915 8142
rect 475 7147 1690 7148
rect 398 7131 1690 7147
rect 398 6950 411 7131
rect 572 7124 1690 7131
rect 572 6950 1249 7124
rect 398 1040 424 6950
rect 491 6941 1249 6950
rect 1662 6941 1690 7124
rect 491 6924 1690 6941
rect 491 1040 505 6924
rect 1844 6839 1915 7884
rect 1619 6837 2084 6839
rect 640 6817 2084 6837
rect 640 6766 1648 6817
rect 572 6626 1231 6688
rect 655 6276 800 6551
rect 655 6263 994 6276
rect 559 6202 603 6251
rect 1087 6202 1131 6253
rect 559 6140 1131 6202
rect 559 6097 603 6140
rect 559 4297 603 5761
rect 651 4123 812 6085
rect 879 4039 1039 5816
rect 1087 4039 1131 6140
rect 643 4002 1131 4039
rect 879 3980 1039 4002
rect 556 3795 602 3973
rect 556 3787 1042 3795
rect 1084 3787 1130 3972
rect 1183 3787 1231 6626
rect 1619 6446 1648 6766
rect 2061 6446 2084 6817
rect 1619 6421 2084 6446
rect 2153 6188 2186 10082
rect 1842 6130 2186 6188
rect 2244 6188 2365 10082
rect 2447 6188 2499 6189
rect 2244 6130 2499 6188
rect 1842 5292 1991 6130
rect 1842 4345 1865 5292
rect 556 3713 1610 3787
rect 649 3511 1410 3570
rect 649 3500 1048 3511
rect 562 3374 1231 3447
rect 880 3007 1026 3314
rect 555 2958 599 3004
rect 1087 2958 1128 3004
rect 555 2936 1128 2958
rect 555 2880 1131 2936
rect 555 2843 599 2880
rect 398 638 505 1040
rect 555 832 599 2512
rect 540 815 602 832
rect 540 723 602 733
rect 656 641 792 2835
rect 398 183 415 638
rect 483 183 505 638
rect 896 581 1031 2551
rect 1087 832 1131 2880
rect 1078 815 1140 832
rect 1078 723 1140 733
rect 1087 581 1131 723
rect 644 535 1131 581
rect 896 516 1031 535
rect 574 390 1116 450
rect 557 389 1116 390
rect 557 296 646 389
rect 1043 327 1130 389
rect 660 296 1130 327
rect 1183 296 1231 3374
rect 1340 2466 1410 3511
rect 1519 2856 1610 3713
rect 1842 3234 1991 4345
rect 2431 3234 2499 6130
rect 1842 3181 2499 3234
rect 2358 2965 2499 3181
rect 1519 2781 2111 2856
rect 1735 2770 2111 2781
rect 1637 2707 1681 2752
rect 2151 2707 2195 2753
rect 1637 2643 2195 2707
rect 1637 2466 1681 2643
rect 2151 2599 2195 2643
rect 1340 2396 1869 2466
rect 1610 2365 1681 2396
rect 1610 2279 1681 2289
rect 1637 795 1681 2279
rect 1732 735 1869 2396
rect 1939 648 2105 2574
rect 2151 2364 2224 2374
rect 2151 2279 2224 2289
rect 2151 795 2195 2279
rect 2358 648 2364 2965
rect 1712 519 2364 648
rect 2493 519 2499 2965
rect 2658 2854 2868 2867
rect 2658 2662 2669 2854
rect 2855 2662 2868 2854
rect 2658 2649 2868 2662
rect 1712 477 2115 519
rect 2358 507 2499 519
rect 2740 413 2794 2649
rect 1651 359 2794 413
rect 2358 300 2499 315
rect 557 277 1563 296
rect 1715 277 2111 296
rect 557 232 2111 277
rect 1436 199 2111 232
rect 398 71 409 183
rect 494 71 505 183
rect 398 54 505 71
rect 2358 62 2366 300
rect 2492 147 2499 300
rect 3336 147 3936 10819
rect 4336 147 4936 10819
rect 5336 147 5936 10819
rect 6336 147 6936 10819
rect 7336 147 7936 10819
rect 8585 147 8673 10819
rect 2492 62 8673 147
rect 0 0 140 40
rect 2358 39 8673 62
<< via1 >>
rect 44 106 116 11762
rect 432 7332 531 10816
rect 956 10833 1010 10919
rect 956 10799 1001 10833
rect 1001 10799 1010 10833
rect 956 10767 1010 10799
rect 631 10152 685 10304
rect 877 8353 936 8533
rect 1141 8632 1235 10663
rect 1141 7320 1235 8357
rect 1396 11256 1437 11802
rect 1437 11256 1556 11802
rect 1608 11731 4718 11802
rect 5004 11731 8605 11802
rect 2645 11482 4893 11550
rect 4950 11498 8431 11566
rect 1797 11363 2413 11379
rect 1797 11323 1814 11363
rect 1814 11323 2405 11363
rect 2405 11323 2413 11363
rect 1797 11310 2413 11323
rect 2014 11031 8634 11105
rect 1385 8616 1560 10764
rect 1850 10521 1919 10686
rect 2177 10545 2248 10923
rect 2424 10247 2497 10714
rect 1806 8453 2000 8520
rect 1385 7185 1560 8334
rect 424 6950 491 7107
rect 424 1040 491 6950
rect 1648 6446 2061 6817
rect 2186 6130 2244 10082
rect 2186 5438 2244 6130
rect 1865 4345 1991 5292
rect 1991 4345 2414 5292
rect 540 733 602 815
rect 415 183 483 638
rect 1078 733 1140 815
rect 1610 2289 1681 2365
rect 2151 2289 2224 2364
rect 415 74 483 183
<< metal2 >>
rect 0 11762 140 11832
rect 0 106 44 11762
rect 116 106 140 11762
rect 406 10816 559 10855
rect 406 7332 432 10816
rect 531 7332 559 10816
rect 768 10445 828 11911
rect 943 10767 956 10919
rect 1010 10866 1023 10919
rect 1133 10866 1193 11912
rect 1010 10806 1193 10866
rect 1360 11802 4740 11840
rect 1360 11256 1396 11802
rect 1556 11731 1608 11802
rect 4718 11731 4740 11802
rect 1556 11689 4740 11731
rect 1556 11256 1590 11689
rect 4816 11591 4917 11911
rect 4978 11802 8641 11840
rect 4978 11731 5004 11802
rect 8605 11731 8641 11802
rect 4978 11689 8641 11731
rect 4816 11582 8453 11591
rect 2619 11566 8453 11582
rect 2619 11550 4950 11566
rect 2619 11482 2645 11550
rect 4893 11498 4950 11550
rect 8431 11498 8453 11566
rect 4893 11482 8453 11498
rect 2619 11481 8453 11482
rect 2619 11460 4916 11481
rect 1782 11379 2440 11386
rect 1782 11310 1797 11379
rect 2413 11310 2440 11379
rect 1782 11304 2440 11310
rect 1010 10767 1023 10806
rect 1360 10764 1590 11256
rect 618 10385 828 10445
rect 1114 10663 1267 10681
rect 618 10304 698 10385
rect 618 10152 631 10304
rect 685 10152 698 10304
rect 618 10144 698 10152
rect 1114 8632 1141 10663
rect 1235 8632 1267 10663
rect 1114 8602 1267 8632
rect 1360 8616 1385 10764
rect 1560 10445 1590 10764
rect 1850 10686 1919 11304
rect 1968 11105 8670 11128
rect 1968 11031 2014 11105
rect 8634 11031 8670 11105
rect 1968 10980 8670 11031
rect 1850 10512 1919 10521
rect 2153 10923 2366 10980
rect 2153 10545 2177 10923
rect 2248 10545 2366 10923
rect 2153 10508 2366 10545
rect 2414 10714 2508 10730
rect 2414 10445 2424 10714
rect 1560 10247 2424 10445
rect 2497 10247 2508 10714
rect 1560 10235 2508 10247
rect 1560 8616 1590 10235
rect 1141 8601 1235 8602
rect 1360 8581 1590 8616
rect 2161 10082 2359 10130
rect 867 8353 877 8533
rect 936 8514 946 8533
rect 1796 8514 1806 8520
rect 936 8457 1806 8514
rect 936 8353 946 8457
rect 1796 8453 1806 8457
rect 2000 8453 2010 8520
rect 1114 8357 1267 8388
rect 406 7298 559 7332
rect 1114 7320 1141 8357
rect 1235 7320 1267 8357
rect 1114 7293 1267 7320
rect 1360 8334 1590 8369
rect 1360 7185 1385 8334
rect 1560 7185 1590 8334
rect 1360 7155 1590 7185
rect 397 7107 624 7146
rect 397 7105 424 7107
rect 491 7105 624 7107
rect 397 999 423 7105
rect 0 0 140 106
rect 398 900 423 999
rect 580 900 624 7105
rect 1619 6817 2084 6839
rect 1619 6446 1648 6817
rect 2061 6446 2084 6817
rect 1619 6421 2084 6446
rect 2161 5438 2186 10082
rect 2244 5438 2359 10082
rect 2161 5312 2359 5438
rect 1816 5292 2435 5312
rect 1816 4345 1835 5292
rect 2414 4345 2435 5292
rect 1816 4322 2435 4345
rect 1600 2289 1610 2365
rect 1681 2354 1691 2365
rect 2141 2354 2151 2364
rect 1681 2302 2151 2354
rect 1681 2289 1691 2302
rect 2141 2289 2151 2302
rect 2224 2289 2234 2364
rect 398 880 624 900
rect 398 668 497 880
rect 530 733 540 815
rect 602 799 612 815
rect 1068 799 1078 815
rect 602 743 1078 799
rect 602 733 612 743
rect 1068 733 1078 743
rect 1140 733 1150 815
rect 398 648 623 668
rect 398 638 423 648
rect 398 74 415 638
rect 580 91 623 648
rect 483 74 623 91
rect 398 52 623 74
<< via2 >>
rect 44 106 116 11762
rect 432 7332 531 10816
rect 1141 8632 1235 10663
rect 1141 7320 1235 8357
rect 423 1040 424 7105
rect 424 1040 491 7105
rect 491 1040 580 7105
rect 423 900 580 1040
rect 1648 6446 2061 6817
rect 1835 4345 1865 5292
rect 1865 4345 2162 5292
rect 423 638 580 648
rect 423 91 483 638
rect 483 91 580 638
<< metal3 >>
rect 0 11762 246 11911
rect 0 11727 44 11762
rect 116 11727 246 11762
rect 0 93 10 11727
rect 130 93 246 11727
rect 406 10816 559 10855
rect 406 7332 432 10816
rect 531 7332 559 10816
rect 406 7298 559 7332
rect 1114 10663 1267 10681
rect 1114 7320 1141 10663
rect 1235 7320 1267 10663
rect 1114 7293 1267 7320
rect 0 0 246 93
rect 401 7105 719 7140
rect 401 900 423 7105
rect 580 7087 719 7105
rect 401 648 440 900
rect 401 91 423 648
rect 401 87 440 91
rect 684 87 719 7087
rect 1619 6817 2084 6839
rect 1619 6446 1648 6817
rect 2061 6446 2084 6817
rect 1619 6422 2084 6446
rect 1367 5292 2190 5313
rect 1367 5282 1835 5292
rect 1367 4364 1407 5282
rect 1367 4345 1835 4364
rect 2162 4345 2190 5292
rect 1367 4321 2190 4345
rect 1367 4125 2433 4321
rect 401 52 719 87
<< via3 >>
rect 10 106 44 11727
rect 44 106 116 11727
rect 116 106 130 11727
rect 10 93 130 106
rect 432 7942 531 10816
rect 1141 8632 1235 10663
rect 1141 8357 1235 8632
rect 1141 7320 1235 8357
rect 440 900 580 7087
rect 580 900 684 7087
rect 440 648 684 900
rect 440 91 580 648
rect 580 91 684 648
rect 440 87 684 91
rect 1648 6446 2061 6817
rect 1407 4364 1835 5282
rect 1835 4364 2126 5282
<< metal4 >>
rect 0 11727 246 11911
rect 0 93 10 11727
rect 130 7750 246 11727
rect 393 10816 722 11911
rect 910 11160 2093 11192
rect 910 10893 929 11160
rect 2069 10893 2093 11160
rect 910 10857 2093 10893
rect 393 7942 432 10816
rect 531 7942 722 10816
rect 393 7932 722 7942
rect 1029 10663 1429 10681
rect 1029 7750 1141 10663
rect 130 7320 1141 7750
rect 1235 7320 1429 10663
rect 130 7262 1429 7320
rect 130 93 246 7262
rect 0 0 246 93
rect 401 7087 719 7140
rect 401 87 440 7087
rect 684 87 719 7087
rect 401 0 719 87
rect 1029 5313 1429 6998
rect 1610 6817 2093 10857
rect 1610 6446 1648 6817
rect 2061 6446 2093 6817
rect 1610 6400 2093 6446
rect 1029 5282 2162 5313
rect 1029 4364 1407 5282
rect 2126 4364 2162 5282
rect 1029 4025 2162 4364
rect 2433 4115 8633 4807
rect 1029 3831 8633 4025
rect 1029 0 1429 3831
<< via4 >>
rect 929 10893 2069 11160
rect 1437 4364 2126 5282
<< metal5 >>
rect 905 11160 2442 11185
rect 905 10893 929 11160
rect 2069 10893 2442 11160
rect 905 10865 2442 10893
rect 1367 5282 2549 5313
rect 1367 4364 1437 5282
rect 2126 4521 2549 5282
rect 2126 4364 2190 4521
rect 1367 4327 2190 4364
use sky130_fd_pr__cap_mim_m3_1_WRT4AW  sky130_fd_pr__cap_mim_m3_1_WRT4AW_0 primitives
timestamp 1606502073
transform 0 -1 5533 -1 0 7041
box -3136 -3100 3136 3100
use sky130_fd_pr__cap_mim_m3_2_W5U4AW  sky130_fd_pr__cap_mim_m3_2_W5U4AW_0 primitives
timestamp 1606502073
transform 0 -1 5533 1 0 7984
box -3179 -3101 3201 3101
use sky130_fd_pr__nfet_g5v0d10v5_PKVMTM  sky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0 primitives
timestamp 1625577137
transform 0 -1 1914 1 0 2674
box -308 -458 308 458
use sky130_fd_pr__nfet_g5v0d10v5_TGFUGS  sky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 primitives
timestamp 1606063140
transform 0 -1 1915 1 0 1529
box -962 -458 962 458
use sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC  sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1 primitives
timestamp 1605994897
transform 0 -1 1915 -1 0 385
box -308 -458 308 458
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0 primitives
timestamp 1606063140
transform 0 -1 843 1 0 3406
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1
timestamp 1606063140
transform 0 -1 843 1 0 3892
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2
timestamp 1606063140
transform 0 -1 843 1 0 6658
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3
timestamp 1606063140
transform 0 -1 843 1 0 422
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YEUEBV  sky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 primitives
timestamp 1606063140
transform 0 -1 843 1 0 5032
box -992 -497 992 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPBG  sky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 primitives
timestamp 1606063140
transform 0 -1 843 1 0 2920
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPXE  sky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 primitives
timestamp 1606063140
transform 0 -1 843 1 0 6172
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ  sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 primitives
timestamp 1606063140
transform 0 -1 843 1 0 1671
box -1101 -497 1101 497
use sky130_fd_pr__res_xhigh_po_0p69_S5N9F3  sky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0 primitives
timestamp 1606074388
transform 0 -1 5586 1 0 5460
box -5446 -3098 5446 3098
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 -1 2280 1 0 8537
box -66 -43 1986 897
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_1
timestamp 1746753973
transform 0 -1 1246 1 0 7491
box -66 -43 1986 897
use sky130_fd_sc_hvl__buf_32  sky130_fd_sc_hvl__buf_32_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 1 0 1539 0 1 11003
box -66 -43 6786 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 1 0 8259 0 1 11003
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_1
timestamp 1746753973
transform 0 -1 2280 -1 0 10841
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_2
timestamp 1746753973
transform 0 -1 1246 -1 0 11235
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_3
timestamp 1746753973
transform 0 -1 1246 -1 0 11619
box -66 -43 450 897
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 -1 1246 1 0 9411
box -66 -43 1506 897
use sky130_fd_sc_hvl__schmittbuf_1  sky130_fd_sc_hvl__schmittbuf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 -1 2280 1 0 7481
box -66 -43 1122 897
<< labels >>
flabel metal4 s 401 0 719 7140 0 FreeSans 320 270 0 0 vdd3v3
port 0 nsew power bidirectional
flabel metal4 s 393 7932 722 11912 0 FreeSans 320 270 0 0 vdd1v8
port 1 nsew power bidirectional
flabel metal4 s 0 0 246 11911 0 FreeSans 800 270 0 0 vss1v8
port 7 nsew ground bidirectional
flabel metal4 s 1029 0 1429 6998 0 FreeSans 320 270 0 0 vss3v3
port 2 nsew ground bidirectional
flabel metal2 1133 11723 1193 11912 0 FreeSans 320 270 0 0 por_l
port 5 nsew signal output
flabel metal2 768 11722 828 11911 0 FreeSans 320 270 0 0 porb_l
port 6 nsew signal output
flabel metal2 4816 11574 4917 11911 0 FreeSans 320 270 0 0 porb_h
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 8715 11912
string LEFclass BLOCK
string MASKHINTS_HVI 300 7390 2370 11900 2370 10915 8755 11900
<< end >>
