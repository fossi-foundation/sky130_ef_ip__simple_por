VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__simple_por
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__simple_por ;
  ORIGIN 0.000 0.000 ;
  SIZE 63.720 BY 41.690 ;
  PIN vdd3v3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.190 39.825 0.365 41.415 ;
    END
  END vdd3v3
  PIN vdd1v8
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 54.010 39.810 55.900 41.455 ;
    END
  END vdd1v8
  PIN vss3v3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.190 36.275 21.750 38.275 ;
    END
  END vss3v3
  PIN porb_h
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 54.545 33.825 56.710 34.170 ;
    END
  END porb_h
  PIN por_l
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 53.960 37.455 56.720 37.755 ;
    END
  END por_l
  PIN porb_l
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 51.855 39.280 56.715 39.580 ;
    END
  END porb_l
  PIN vss1v8
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.070 42.720 0.290 43.420 ;
    END
  END vss1v8
  OBS
      LAYER li1 ;
        RECT -0.070 42.760 56.090 43.380 ;
        RECT 0.000 0.180 56.090 41.690 ;
      LAYER met1 ;
        RECT 0.290 42.720 56.090 43.420 ;
        RECT 0.125 0.055 56.090 41.690 ;
      LAYER met2 ;
        RECT -0.070 42.720 56.090 43.420 ;
        RECT 0.000 30.880 56.090 41.690 ;
      LAYER met3 ;
        RECT -0.070 42.190 56.070 43.420 ;
        RECT 0.000 39.980 56.070 41.690 ;
        RECT 0.000 38.880 51.455 39.980 ;
        RECT 0.000 38.155 56.070 38.880 ;
        RECT 0.000 37.055 53.560 38.155 ;
        RECT 0.000 34.570 56.070 37.055 ;
        RECT 0.000 33.425 54.145 34.570 ;
        RECT 0.000 0.255 56.070 33.425 ;
      LAYER met4 ;
        RECT 36.240 41.690 38.680 43.420 ;
        RECT 0.765 39.425 53.610 41.690 ;
        RECT 0.365 39.410 53.610 39.425 ;
        RECT 0.365 38.675 55.890 39.410 ;
        RECT 22.150 35.875 55.890 38.675 ;
        RECT 0.365 0.255 55.890 35.875 ;
      LAYER met5 ;
        RECT 21.565 0.250 55.855 38.895 ;
  END
END sky130_ef_ip__simple_por
END LIBRARY

