magic
tech sky130A
magscale 1 2
timestamp 1638030790
<< obsli1 >>
rect -14 8552 11218 8676
rect 0 36 11218 8338
<< metal1 >>
rect -14 8544 58 8684
<< obsm1 >>
rect 58 8544 11218 8684
rect 25 11 11218 8338
<< obsm2 >>
rect 38 6176 10918 8287
<< metal3 >>
rect 10371 7856 11343 7916
rect 10792 7491 11344 7551
rect 10909 6765 11342 6834
<< obsm3 >>
rect 38 7996 10918 8283
rect 38 7776 10291 7996
rect 38 7631 10918 7776
rect 38 7411 10712 7631
rect 38 6914 10918 7411
rect 38 6685 10829 6914
rect 38 51 10918 6685
<< metal4 >>
rect 38 7965 7241 8283
rect 7356 7962 11180 8291
rect 38 7255 4350 7655
<< obsm4 >>
rect 73 7882 4430 7885
rect 73 7735 11178 7882
rect 4430 7175 11178 7735
rect 73 51 11178 7175
<< obsm5 >>
rect 4313 50 11171 7779
<< labels >>
rlabel metal4 s 38 7255 4350 7655 6 vss3v3
port 3 nsew ground bidirectional
rlabel metal3 s 10909 6765 11342 6834 6 porb_h
port 4 nsew signal output
rlabel metal3 s 10792 7491 11344 7551 6 por_l
port 5 nsew signal output
rlabel metal3 s 10371 7856 11343 7916 6 porb_l
port 6 nsew signal output
rlabel metal1 s -14 8544 58 8684 6 vss1v8
port 7 nsew ground bidirectional
rlabel metal4 7356 7962 11180 8291 0 vdd1v8
port 1 nsew power bidirectional
rlabel metal4 38 7965 7241 8283 0 vdd3v3
port 2 nsew power bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 11344 8338
string GDS_FILE ../gds/sky130_ef_ip__simple_por.gds
string GDS_START 0
string LEFview TRUE
<< end >>
